module RAMB36E2 (
  CASDOUTA,
  CASDOUTB,
  CASDOUTPA,
  CASDOUTPB,
  CASOUTDBITERR,
  CASOUTSBITERR,
  DBITERR,
  DOUTADOUT,
  DOUTBDOUT,
  DOUTPADOUTP,
  DOUTPBDOUTP,
  ECCPARITY,
  RDADDRECC,
  SBITERR,

  ADDRARDADDR,
  ADDRBWRADDR,
  ADDRENA,
  ADDRENB,
  CASDIMUXA,
  CASDIMUXB,
  CASDINA,
  CASDINB,
  CASDINPA,
  CASDINPB,
  CASDOMUXA,
  CASDOMUXB,
  CASDOMUXEN_A,
  CASDOMUXEN_B,
  CASINDBITERR,
  CASINSBITERR,
  CASOREGIMUXA,
  CASOREGIMUXB,
  CASOREGIMUXEN_A,
  CASOREGIMUXEN_B,
  CLKARDCLK,
  CLKBWRCLK,
  DINADIN,
  DINBDIN,
  DINPADINP,
  DINPBDINP,
  ECCPIPECE,
  ENARDEN,
  ENBWREN,
  INJECTDBITERR,
  INJECTSBITERR,
  REGCEAREGCE,
  REGCEB,
  RSTRAMARSTRAM,
  RSTRAMB,
  RSTREGARSTREG,
  RSTREGB,
  SLEEP,
  WEA,
  WEBWE
);

  parameter CASCADE_ORDER_A = "NONE";
  parameter CASCADE_ORDER_B = "NONE";
  parameter CLOCK_DOMAINS = "INDEPENDENT";
  parameter integer DOA_REG = 1;
  parameter integer DOB_REG = 1;
  parameter ENADDRENA = "FALSE";
  parameter ENADDRENB = "FALSE";
  parameter EN_ECC_PIPE = "FALSE";
  parameter EN_ECC_READ = "FALSE";
  parameter EN_ECC_WRITE = "FALSE";
  parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [35:0] INIT_A = 36'h000000000;
  parameter [35:0] INIT_B = 36'h000000000;
  parameter INIT_FILE = "NONE";
  parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
  parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
  parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
  parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
  parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
  parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
  parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
  parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
  parameter RDADDRCHANGEA = "FALSE";
  parameter RDADDRCHANGEB = "FALSE";
  parameter integer READ_WIDTH_A = 0;
  parameter integer READ_WIDTH_B = 0;
  parameter RSTREG_PRIORITY_A = "RSTREG";
  parameter RSTREG_PRIORITY_B = "RSTREG";
  parameter SIM_COLLISION_CHECK = "ALL";
  parameter SLEEP_ASYNC = "FALSE";
  parameter [35:0] SRVAL_A = 36'h000000000;
  parameter [35:0] SRVAL_B = 36'h000000000;
  parameter WRITE_MODE_A = "NO_CHANGE";
  parameter WRITE_MODE_B = "NO_CHANGE";
  parameter integer WRITE_WIDTH_A = 0;
  parameter integer WRITE_WIDTH_B = 0;
  
  output [31:0] CASDOUTA;
  output [31:0] CASDOUTB;
  output [3:0] CASDOUTPA;
  output [3:0] CASDOUTPB;
  output CASOUTDBITERR;
  output CASOUTSBITERR;
  output DBITERR;
  output [31:0] DOUTADOUT;
  output [31:0] DOUTBDOUT;
  output [3:0] DOUTPADOUTP;
  output [3:0] DOUTPBDOUTP;
  output [7:0] ECCPARITY;
  output [8:0] RDADDRECC;
  output SBITERR;

  input [14:0] ADDRARDADDR;
  input [14:0] ADDRBWRADDR;
  input ADDRENA;
  input ADDRENB;
  input CASDIMUXA;
  input CASDIMUXB;
  input [31:0] CASDINA;
  input [31:0] CASDINB;
  input [3:0] CASDINPA;
  input [3:0] CASDINPB;
  input CASDOMUXA;
  input CASDOMUXB;
  input CASDOMUXEN_A;
  input CASDOMUXEN_B;
  input CASINDBITERR;
  input CASINSBITERR;
  input CASOREGIMUXA;
  input CASOREGIMUXB;
  input CASOREGIMUXEN_A;
  input CASOREGIMUXEN_B;
  input CLKARDCLK;
  input CLKBWRCLK;
  input [31:0] DINADIN;
  input [31:0] DINBDIN;
  input [3:0] DINPADINP;
  input [3:0] DINPBDINP;
  input ECCPIPECE;
  input ENARDEN;
  input ENBWREN;
  input INJECTDBITERR;
  input INJECTSBITERR;
  input REGCEAREGCE;
  input REGCEB;
  input RSTRAMARSTRAM;
  input RSTRAMB;
  input RSTREGARSTREG;
  input RSTREGB;
  input SLEEP;
  input [3:0] WEA;
  input [7:0] WEBWE;
  
  localparam [ 0:0] SYNC_FIFO1_i  = 1'd0;
  localparam [ 0:0] FMODE1_i      = 1'd0;
  localparam [ 0:0] POWERDN1_i    = 1'd0;
  localparam [ 0:0] SLEEP1_i      = 1'd0;
  localparam [ 0:0] PROTECT1_i    = 1'd0;
  localparam [11:0] UPAE1_i       = 12'd10;
  localparam [11:0] UPAF1_i       = 12'd10;
  
  localparam [ 0:0] SYNC_FIFO2_i  = 1'd0;
  localparam [ 0:0] FMODE2_i      = 1'd0;
  localparam [ 0:0] POWERDN2_i    = 1'd0;
  localparam [ 0:0] SLEEP2_i      = 1'd0;
  localparam [ 0:0] PROTECT2_i    = 1'd0;
  localparam [10:0] UPAE2_i       = 11'd10;
  localparam [10:0] UPAF2_i       = 11'd10;
  
  assign CASDOUTA =32'h0;
  assign CASDOUTB =32'h0;
  assign CASDOUTPA =4'h0;
  assign CASDOUTPB =4'h0;
  
  assign CASOUTDBITERR = 1'b0; 
  assign CASOUTSBITERR = 1'b0; 
  assign DBITERR = 1'b0; 
  assign SBITERR = 1'b0; 

  assign ECCPARITY =8'h0;
  assign RDADDRECC =9'h0;

  
  function [2:0] mode;
	input integer width;
	case (width)
		1: mode = 3'b101;
		2: mode = 3'b110;
		4: mode = 3'b100;
		8,9: mode = 3'b001;
		16, 18: mode = 3'b010;
		32, 36: mode = 3'b011;
		default: mode = 3'b000;
	endcase
  endfunction
  
  localparam [ 2:0] RMODE_A1_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] WMODE_A1_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] RMODE_A2_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] WMODE_A2_i    = mode(READ_WIDTH_A);

  localparam [ 2:0] RMODE_B1_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] WMODE_B1_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] RMODE_B2_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] WMODE_B2_i    = mode(WRITE_WIDTH_B);
  
    TDP36K bram32k_0 (
	.RESET_ni(),
	.WEN_A1_i(WEA[0]),
	.WEN_B1_i(WEBWE[0]),
	.REN_A1_i(ENARDEN),
	.REN_B1_i(1'b0),
	.CLK_A1_i(CLKARDCLK),
	.CLK_B1_i(CLKBWRCLK),
	.BE_A1_i({WEA[1:0]}),
	.BE_B1_i({WEBWE[1:0]}),
	.ADDR_A1_i(ADDRARDADDR),
	.ADDR_B1_i(ADDRBWRADDR),
	.WDATA_A1_i({DINPADINP[1:0],DINADIN[15:0]}),
	.WDATA_B1_i({DINPBDINP[1:0],DINBDIN[15:0]}),
	.RDATA_A1_o({DOUTPADOUTP[1:0],DOUTADOUT[15:0]}),
	.RDATA_B1_o({DOUTPBDOUTP[1:0],DOUTBDOUT[15:0]}),
	.FLUSH1_i(1'b0),
	.WEN_A2_i(1'b0),
	.WEN_B2_i(1'b0),
	.REN_A2_i(1'b0),
	.REN_B2_i(1'b0),
	.CLK_A2_i(),
	.CLK_B2_i(),
	.BE_A2_i({WEA[3:2]}),
	.BE_B2_i({WEBWE[3:2]}),
	.ADDR_A2_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.ADDR_B2_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.WDATA_A2_i({DINPADINP[3:2],DINADIN[31:16]}),
	.WDATA_B2_i({DINPBDINP[3:2],DINBDIN[31:16]}),
	.RDATA_A2_o({DOUTPADOUTP[3:2],DOUTADOUT[31:16]}),
	.RDATA_B2_o({DOUTPBDOUTP[3:2],DOUTBDOUT[31:16]}),
	.FLUSH2_i(1'b0)
	);
	defparam bram32k_0.MODE_BITS = { 1'b0,
		UPAF2_i, UPAE2_i, PROTECT2_i, SLEEP2_i, POWERDN2_i, FMODE2_i, WMODE_B2_i, WMODE_A2_i, RMODE_B2_i, RMODE_A2_i, SYNC_FIFO2_i,
		UPAF1_i, UPAE1_i, PROTECT1_i, SLEEP1_i, POWERDN1_i, FMODE1_i, WMODE_B1_i, WMODE_A1_i, RMODE_B1_i, RMODE_A1_i, SYNC_FIFO1_i
	};

endmodule

module RAMB18E2 (
  CASDOUTA,
  CASDOUTB,
  CASDOUTPA,
  CASDOUTPB,
  DOUTADOUT,
  DOUTBDOUT,
  DOUTPADOUTP,
  DOUTPBDOUTP,

  ADDRARDADDR,
  ADDRBWRADDR,
  ADDRENA,
  ADDRENB,
  CASDIMUXA,
  CASDIMUXB,
  CASDINA,
  CASDINB,
  CASDINPA,
  CASDINPB,
  CASDOMUXA,
  CASDOMUXB,
  CASDOMUXEN_A,
  CASDOMUXEN_B,
  CASOREGIMUXA,
  CASOREGIMUXB,
  CASOREGIMUXEN_A,
  CASOREGIMUXEN_B,
  CLKARDCLK,
  CLKBWRCLK,
  DINADIN,
  DINBDIN,
  DINPADINP,
  DINPBDINP,
  ENARDEN,
  ENBWREN,
  REGCEAREGCE,
  REGCEB,
  RSTRAMARSTRAM,
  RSTRAMB,
  RSTREGARSTREG,
  RSTREGB,
  SLEEP,
  WEA,
  WEBWE
);

  parameter CASCADE_ORDER_A = "NONE";
  parameter CASCADE_ORDER_B = "NONE";
  parameter CLOCK_DOMAINS = "INDEPENDENT";
  parameter integer DOA_REG = 1;
  parameter integer DOB_REG = 1;
  parameter ENADDRENA = "FALSE";
  parameter ENADDRENB = "FALSE";
  parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter [17:0] INIT_A = 18'h00000;
  parameter [17:0] INIT_B = 18'h00000;
  parameter INIT_FILE = "NONE";
  parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
  parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
  parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
  parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
  parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
  parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
  parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
  parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
  parameter RDADDRCHANGEA = "FALSE";
  parameter RDADDRCHANGEB = "FALSE";
  parameter integer READ_WIDTH_A = 0;
  parameter integer READ_WIDTH_B = 0;
  parameter RSTREG_PRIORITY_A = "RSTREG";
  parameter RSTREG_PRIORITY_B = "RSTREG";
  parameter SIM_COLLISION_CHECK = "ALL";
  parameter SLEEP_ASYNC = "FALSE";
  parameter [17:0] SRVAL_A = 18'h00000;
  parameter [17:0] SRVAL_B = 18'h00000;
  parameter WRITE_MODE_A = "NO_CHANGE";
  parameter WRITE_MODE_B = "NO_CHANGE";
  parameter integer WRITE_WIDTH_A = 0;
  parameter integer WRITE_WIDTH_B = 0;
  
  output [15:0] CASDOUTA;
  output [15:0] CASDOUTB;
  output [1:0] CASDOUTPA;
  output [1:0] CASDOUTPB;
  output [15:0] DOUTADOUT;
  output [15:0] DOUTBDOUT;
  output [1:0] DOUTPADOUTP;
  output [1:0] DOUTPBDOUTP;

  input [13:0] ADDRARDADDR;
  input [13:0] ADDRBWRADDR;
  input ADDRENA;
  input ADDRENB;
  input CASDIMUXA;
  input CASDIMUXB;
  input [15:0] CASDINA;
  input [15:0] CASDINB;
  input [1:0] CASDINPA;
  input [1:0] CASDINPB;
  input CASDOMUXA;
  input CASDOMUXB;
  input CASDOMUXEN_A;
  input CASDOMUXEN_B;
  input CASOREGIMUXA;
  input CASOREGIMUXB;
  input CASOREGIMUXEN_A;
  input CASOREGIMUXEN_B;
  input CLKARDCLK;
  input CLKBWRCLK;
  input [15:0] DINADIN;
  input [15:0] DINBDIN;
  input [1:0] DINPADINP;
  input [1:0] DINPBDINP;
  input ENARDEN;
  input ENBWREN;
  input REGCEAREGCE;
  input REGCEB;
  input RSTRAMARSTRAM;
  input RSTRAMB;
  input RSTREGARSTREG;
  input RSTREGB;
  input SLEEP;
  input [1:0] WEA;
  input [3:0] WEBWE;
  
  localparam [ 0:0] SYNC_FIFO1_i  = 1'd0;
  localparam [ 0:0] FMODE1_i      = 1'd0;
  localparam [ 0:0] POWERDN1_i    = 1'd0;
  localparam [ 0:0] SLEEP1_i      = 1'd0;
  localparam [ 0:0] PROTECT1_i    = 1'd0;
  localparam [11:0] UPAE1_i       = 12'd10;
  localparam [11:0] UPAF1_i       = 12'd10;
  
  localparam [ 0:0] SYNC_FIFO2_i  = 1'd0;
  localparam [ 0:0] FMODE2_i      = 1'd0;
  localparam [ 0:0] POWERDN2_i    = 1'd0;
  localparam [ 0:0] SLEEP2_i      = 1'd0;
  localparam [ 0:0] PROTECT2_i    = 1'd0;
  localparam [10:0] UPAE2_i       = 11'd10;
  localparam [10:0] UPAF2_i       = 11'd10;
  
  assign CASDOUTA =16'h0;
  assign CASDOUTB =16'h0;
  assign CASDOUTPA =2'h0;
  assign CASDOUTPB =2'h0;
   
  function [2:0] mode;
	input integer width;
	case (width)
		1: mode = 3'b101;
		2: mode = 3'b110;
		4: mode = 3'b100;
		8,9: mode = 3'b001;
		16, 18: mode = 3'b010;
		32, 36: mode = 3'b011;
		default: mode = 3'b000;
	endcase
  endfunction
  
  localparam [ 2:0] RMODE_A1_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] WMODE_A1_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] RMODE_A2_i    = mode(READ_WIDTH_A);
  localparam [ 2:0] WMODE_A2_i    = mode(READ_WIDTH_A);

  localparam [ 2:0] RMODE_B1_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] WMODE_B1_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] RMODE_B2_i    = mode(WRITE_WIDTH_B);
  localparam [ 2:0] WMODE_B2_i    = mode(WRITE_WIDTH_B);
  
    TDP36K bram18k_0 (
	.RESET_ni(),
	.WEN_A1_i(WEA[0]),
	.WEN_B1_i(WEBWE[0]),
	.REN_A1_i(ENARDEN),
	.REN_B1_i(1'b0),
	.CLK_A1_i(CLKARDCLK),
	.CLK_B1_i(CLKBWRCLK),
	.BE_A1_i({WEA[1:0]}),
	.BE_B1_i({WEBWE[1:0]}),
	.ADDR_A1_i(ADDRARDADDR),
	.ADDR_B1_i(ADDRBWRADDR),
	.WDATA_A1_i({DINPADINP[1:0],DINADIN[15:0]}),
	.WDATA_B1_i({DINPBDINP[1:0],DINBDIN[15:0]}),
	.RDATA_A1_o({DOUTPADOUTP[1:0],DOUTADOUT[15:0]}),
	.RDATA_B1_o({DOUTPBDOUTP[1:0],DOUTBDOUT[15:0]}),
	.FLUSH1_i(1'b0),
	.WEN_A2_i(1'b0),
	.WEN_B2_i(1'b0),
	.REN_A2_i(1'b0),
	.REN_B2_i(1'b0),
	.CLK_A2_i(),
	.CLK_B2_i(),
	.BE_A2_i({1'b0, 1'b0}),
	.BE_B2_i({WEBWE[3:2]}),
	.ADDR_A2_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.ADDR_B2_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.WDATA_A2_i(18'h0),
	.WDATA_B2_i(18'h0),
	.RDATA_A2_o(),
	.RDATA_B2_o(),
	.FLUSH2_i(1'b0)
	);

	defparam bram18k_0.MODE_BITS = { 1'b0,
		UPAF2_i, UPAE2_i, PROTECT2_i, SLEEP2_i, POWERDN2_i, FMODE2_i, WMODE_B2_i, WMODE_A2_i, RMODE_B2_i, RMODE_A2_i, SYNC_FIFO2_i,
		UPAF1_i, UPAE1_i, PROTECT1_i, SLEEP1_i, POWERDN1_i, FMODE1_i, WMODE_B1_i, WMODE_A1_i, RMODE_B1_i, RMODE_A1_i, SYNC_FIFO1_i
	};

endmodule